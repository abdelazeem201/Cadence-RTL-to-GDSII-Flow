VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER PWdummy
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.3 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.3 ;" ;
END PWdummy

LAYER Nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.6 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.3 ;" ;
END Nwell

LAYER Oxide
  TYPE MASTERSLICE ;
END Oxide

LAYER Nhvt
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
END Nhvt

LAYER Nimp
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
END Nimp

LAYER Phvt
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
END Phvt

LAYER Pimp
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
  SPACING 0 LAYER Nimp ;
END Pimp

LAYER Nzvt
  TYPE IMPLANT ;
  WIDTH 0.35 ;
  SPACING 0.3 ;
END Nzvt

LAYER Nlvt
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
END Nlvt

LAYER Plvt
  TYPE IMPLANT ;
  WIDTH 0.12 ;
  SPACING 0.12 ;
END Plvt

LAYER SiProt
  TYPE IMPLANT ;
  WIDTH 0.22 ;
  SPACING 0.22 ;
END SiProt

LAYER Poly
  TYPE MASTERSLICE ;
END Poly

LAYER Cont
  TYPE CUT ;
  SPACING 0.06 ;
  SPACING 0.08 ADJACENTCUTS 3 WITHIN 0.1 ;
  WIDTH 0.06 ;
  ENCLOSURE BELOW 0.02 0.03 ;
  ENCLOSURE ABOVE 0 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 10 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 10 ) ( 1 10 ) ) ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.06 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.06 0.06 0.06 0.06 0.06 0.06 
    WIDTH 0.1 0.06 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.75 0.06 0.1 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.06 0.1 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.06 0.1 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.06 0.1 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.045 ;
  DIAGSPACING 0.08 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0736 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.15 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.09 WITHIN 0.025 MINLENGTH 0.06 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 1 20 ) ) ;
    ANTENNACUMROUTINGPLUSCUT ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0214 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.1 ADJACENTCUTS 3 WITHIN 0.11 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.005 0.03 ;
  ENCLOSURE ABOVE 0.005 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.19 ;
  WIDTH 0.08 ;
  OFFSET 0.1 0.095 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.32 0.75 1.5 2.5 3.5 
    WIDTH 0 0.07 0.07 0.07 0.07 0.07 0.07 
    WIDTH 0.1 0.07 0.15 0.15 0.15 0.15 0.15 
    WIDTH 0.75 0.07 0.15 0.25 0.25 0.25 0.25 
    WIDTH 1.5 0.07 0.15 0.25 0.45 0.45 0.45 
    WIDTH 2.5 0.07 0.15 0.25 0.45 0.75 0.75 
    WIDTH 3.5 0.07 0.15 0.25 0.45 0.75 1.25 ;
  MINIMUMCUT 1 WIDTH 0.07 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 WITHIN 0.3 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 3 ;
  MINENCLOSEDAREA 0.055 ;
  DIAGSPACING 0.1 ;
  DIAGMINEDGELENGTH 0.1 ;
  RESISTANCE RPERSQ 0.0214 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.1 WITHIN 0.035 MINLENGTH 0.07 PARALLELEDGE 0.08 WITHIN 0.1 ;" ;
END Metal9

LAYER Via9
  TYPE CUT ;
  SPACING 0.18 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.25 ;
  WIDTH 0.18 ;
  ENCLOSURE BELOW 0.015 0.04 ;
  ENCLOSURE ABOVE 0.03 0.05 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.8 ;
END Via9

LAYER Metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.5 0.19 ;
  WIDTH 0.22 ;
  OFFSET 0.6 0.095 ;
  AREA 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.75 1.5 2.5 3.5 
    WIDTH 0 0.2 0.2 0.2 0.2 0.2 
    WIDTH 0.75 0.2 0.35 0.45 0.75 1.25 
    WIDTH 1.5 0.2 0.35 0.45 0.45 0.45 
    WIDTH 2.5 0.2 0.35 0.45 0.75 0.75 
    WIDTH 3.5 0.2 0.35 0.45 0.75 1.25 ;
  MINENCLOSEDAREA 0.11 ;
  RESISTANCE RPERSQ 0.0214 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 8 ;
END Metal10

LAYER Via10
  TYPE CUT ;
  SPACING 0.18 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.25 ;
  WIDTH 0.18 ;
  ENCLOSURE BELOW 0.015 0.04 ;
  ENCLOSURE ABOVE 0.03 0.05 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNACUMAREARATIO 180 ;
  DCCURRENTDENSITY AVERAGE 0.8 ;
END Via10

LAYER Metal11
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.5 0.475 ;
  WIDTH 0.22 ;
  OFFSET 0.6 0.57 ;
  AREA 0.1 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.75 1.5 2.5 3.5 
    WIDTH 0 0.2 0.2 0.2 0.2 0.2 
    WIDTH 0.75 0.2 0.35 0.45 0.75 1.25 
    WIDTH 1.5 0.2 0.35 0.45 0.45 0.45 
    WIDTH 2.5 0.2 0.35 0.45 0.75 0.75 
    WIDTH 3.5 0.2 0.35 0.45 0.75 1.25 ;
  MINENCLOSEDAREA 0.11 ;
  RESISTANCE RPERSQ 0.021 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.099 5000 ) ( 0.1 48045 ) ( 1 48450 ) ) ;
  DCCURRENTDENSITY AVERAGE 8 ;
END Metal11

LAYER Bondpad
  TYPE CUT ;
  PROPERTY LEF58_TYPE "TYPE PASSIVATION ;" ;
  SPACING 8 ;
  WIDTH 55 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 180 ;
END Bondpad

MAXVIASTACK 4 RANGE Metal1 Metal9 ;
VIARULE M11_M10 GENERATE
  LAYER Metal10 ;
    ENCLOSURE 0.015 0.04 ;
  LAYER Metal11 ;
    ENCLOSURE 0.03 0.05 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    SPACING 0.36 BY 0.36 ;
    RESISTANCE 0.040000 ;
END M11_M10

VIARULE M10_M9 GENERATE
  LAYER Metal9 ;
    ENCLOSURE 0.015 0.04 ;
  LAYER Metal10 ;
    ENCLOSURE 0.03 0.05 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    SPACING 0.36 BY 0.36 ;
    RESISTANCE 0.200000 ;
END M10_M9

VIARULE M9_M8 GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal9 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 0.200000 ;
END M9_M8

VIARULE M8_M7 GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M8_M7

VIARULE M7_M6 GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M7_M6

VIARULE M6_M5 GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M6_M5

VIARULE M5_M4 GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M5_M4

VIARULE M4_M3 GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.000000 ;
END M2_M1

VIARULE M1_PO GENERATE
  LAYER Poly ;
    ENCLOSURE 0.02 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 41.000000 ;
END M1_PO

VIARULE M1_DIFF GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.03 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 56.000000 ;
END M1_DIFF

VIARULE M1_PSUB GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.03 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 56.000000 ;
END M1_PSUB

VIARULE M1_PIMP GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.03 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 56.000000 ;
END M1_PIMP

VIARULE M1_NIMP GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.03 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 56.000000 ;
END M1_NIMP

VIARULE M1_NWELL GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.03 0.03 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.03 ;
  LAYER Cont ;
    RECT -0.03 -0.03 0.03 0.03 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 56.000000 ;
END M1_NWELL

VIA M2_M1_HV DEFAULT
  LAYER Metal1 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_HV

VIA M2_M1_VV DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_VV

VIA M2_M1_VH DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal2 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_VH

VIA M2_M1_HH DEFAULT
  LAYER Metal1 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal2 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_HH

VIA M2_M1_2x1_HV_E DEFAULT
  LAYER Metal1 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M2_M1_2x1_HV_E

VIA M2_M1_2x1_HV_W DEFAULT
  LAYER Metal1 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Metal2 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Via1 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_2x1_HV_W

VIA M2_M1_1x2_HV_N DEFAULT
  LAYER Metal1 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M2_M1_1x2_HV_N

VIA M2_M1_1x2_HV_S DEFAULT
  LAYER Metal1 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Metal2 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Via1 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M2_M1_1x2_HV_S

VIA M3_M2_VH DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_VH

VIA M3_M2_HH DEFAULT
  LAYER Metal2 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_HH

VIA M3_M2_HV DEFAULT
  LAYER Metal2 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal3 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_HV

VIA M3_M2_VV DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal3 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_VV

VIA M3_M2_M_NH DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.185 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_M_NH

VIA M3_M2_M_SH DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.185 0.04 0.065 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_M_SH

VIA M3_M2_2x1_VH_E DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M3_M2_2x1_VH_E

VIA M3_M2_2x1_VH_W DEFAULT
  LAYER Metal2 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Metal3 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_2x1_VH_W

VIA M3_M2_1x2_VH_N DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M3_M2_1x2_VH_N

VIA M3_M2_1x2_VH_S DEFAULT
  LAYER Metal2 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Metal3 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Via2 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M3_M2_1x2_VH_S

VIA M4_M3_HV DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_HV

VIA M4_M3_VV DEFAULT
  LAYER Metal3 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_VV

VIA M4_M3_VH DEFAULT
  LAYER Metal3 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal4 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_VH

VIA M4_M3_HH DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal4 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_HH

VIA M4_M3_M_EV DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.185 0.04 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_M_EV

VIA M4_M3_M_WV DEFAULT
  LAYER Metal3 ;
    RECT -0.185 -0.04 0.065 0.04 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_M_WV

VIA M4_M3_2x1_HV_E DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M4_M3_2x1_HV_E

VIA M4_M3_2x1_HV_W DEFAULT
  LAYER Metal3 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Metal4 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_2x1_HV_W

VIA M4_M3_1x2_HV_N DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M4_M3_1x2_HV_N

VIA M4_M3_1x2_HV_S DEFAULT
  LAYER Metal3 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Metal4 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Via3 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M4_M3_1x2_HV_S

VIA M5_M4_VH DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_VH

VIA M5_M4_HH DEFAULT
  LAYER Metal4 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_HH

VIA M5_M4_HV DEFAULT
  LAYER Metal4 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal5 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_HV

VIA M5_M4_VV DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal5 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_VV

VIA M5_M4_M_NH DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.185 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_M_NH

VIA M5_M4_M_SH DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.185 0.04 0.065 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_M_SH

VIA M5_M4_2x1_VH_E DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M5_M4_2x1_VH_E

VIA M5_M4_2x1_VH_W DEFAULT
  LAYER Metal4 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Metal5 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_2x1_VH_W

VIA M5_M4_1x2_VH_N DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Via4 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M5_M4_1x2_VH_N

VIA M5_M4_1x2_VH_S DEFAULT
  LAYER Metal4 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Metal5 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Via4 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M5_M4_1x2_VH_S

VIA M6_M5_HV DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_HV

VIA M6_M5_VV DEFAULT
  LAYER Metal5 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_VV

VIA M6_M5_VH DEFAULT
  LAYER Metal5 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal6 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_VH

VIA M6_M5_HH DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal6 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_HH

VIA M6_M5_M_EV DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.185 0.04 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_M_EV

VIA M6_M5_M_WV DEFAULT
  LAYER Metal5 ;
    RECT -0.185 -0.04 0.065 0.04 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_M_WV

VIA M6_M5_2x1_HV_E DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M6_M5_2x1_HV_E

VIA M6_M5_2x1_HV_W DEFAULT
  LAYER Metal5 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Metal6 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_2x1_HV_W

VIA M6_M5_1x2_HV_N DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Via5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M6_M5_1x2_HV_N

VIA M6_M5_1x2_HV_S DEFAULT
  LAYER Metal5 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Metal6 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Via5 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M6_M5_1x2_HV_S

VIA M7_M6_VH DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_VH

VIA M7_M6_HH DEFAULT
  LAYER Metal6 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_HH

VIA M7_M6_HV DEFAULT
  LAYER Metal6 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal7 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_HV

VIA M7_M6_VV DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal7 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_VV

VIA M7_M6_M_NH DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.185 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_M_NH

VIA M7_M6_M_SH DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.185 0.04 0.065 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_M_SH

VIA M7_M6_2x1_VH_E DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M7_M6_2x1_VH_E

VIA M7_M6_2x1_VH_W DEFAULT
  LAYER Metal6 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Metal7 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_2x1_VH_W

VIA M7_M6_1x2_VH_N DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M7_M6_1x2_VH_N

VIA M7_M6_1x2_VH_S DEFAULT
  LAYER Metal6 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Metal7 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Via6 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M7_M6_1x2_VH_S

VIA M8_M7_HV DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_HV

VIA M8_M7_VV DEFAULT
  LAYER Metal7 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_VV

VIA M8_M7_VH DEFAULT
  LAYER Metal7 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal8 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_VH

VIA M8_M7_HH DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal8 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_HH

VIA M8_M7_M_EV DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.185 0.04 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_M_EV

VIA M8_M7_M_WV DEFAULT
  LAYER Metal7 ;
    RECT -0.185 -0.04 0.065 0.04 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_M_WV

VIA M8_M7_2x1_HV_E DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M8_M7_2x1_HV_E

VIA M8_M7_2x1_HV_W DEFAULT
  LAYER Metal7 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Metal8 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_2x1_HV_W

VIA M8_M7_1x2_HV_N DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M8_M7_1x2_HV_N

VIA M8_M7_1x2_HV_S DEFAULT
  LAYER Metal7 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Metal8 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Via7 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M8_M7_1x2_HV_S

VIA M9_M8_VH DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_VH

VIA M9_M8_HH DEFAULT
  LAYER Metal8 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_HH

VIA M9_M8_HV DEFAULT
  LAYER Metal8 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Metal9 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_HV

VIA M9_M8_VV DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Metal9 ;
    RECT -0.04 -0.065 0.04 0.065 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_VV

VIA M9_M8_M_NH DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.185 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_M_NH

VIA M9_M8_M_SH DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.185 0.04 0.065 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_M_SH

VIA M9_M8_2x1_VH_E DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.18 0.065 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.205 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT 0.105 -0.035 0.175 0.035 ;
END M9_M8_2x1_VH_E

VIA M9_M8_2x1_VH_W DEFAULT
  LAYER Metal8 ;
    RECT -0.18 -0.065 0.04 0.065 ;
  LAYER Metal9 ;
    RECT -0.205 -0.04 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.175 -0.035 -0.105 0.035 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_2x1_VH_W

VIA M9_M8_1x2_VH_N DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.065 0.04 0.205 ;
  LAYER Metal9 ;
    RECT -0.065 -0.04 0.065 0.18 ;
  LAYER Via8 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    RECT -0.035 0.105 0.035 0.175 ;
END M9_M8_1x2_VH_N

VIA M9_M8_1x2_VH_S DEFAULT
  LAYER Metal8 ;
    RECT -0.04 -0.205 0.04 0.065 ;
  LAYER Metal9 ;
    RECT -0.065 -0.18 0.065 0.04 ;
  LAYER Via8 ;
    RECT -0.035 -0.175 0.035 -0.105 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END M9_M8_1x2_VH_S

VIA M10_M9_HV DEFAULT
  LAYER Metal9 ;
    RECT -0.13 -0.105 0.13 0.105 ;
  LAYER Metal10 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_HV

VIA M10_M9_VV DEFAULT
  LAYER Metal9 ;
    RECT -0.105 -0.13 0.105 0.13 ;
  LAYER Metal10 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_VV

VIA M10_M9_VH DEFAULT
  LAYER Metal9 ;
    RECT -0.105 -0.13 0.105 0.13 ;
  LAYER Metal10 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_VH

VIA M10_M9_HH DEFAULT
  LAYER Metal9 ;
    RECT -0.13 -0.105 0.13 0.105 ;
  LAYER Metal10 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_HH

VIA M10_M9_2x1_HV_E DEFAULT
  LAYER Metal9 ;
    RECT -0.13 -0.105 0.49 0.105 ;
  LAYER Metal10 ;
    RECT -0.12 -0.14 0.48 0.14 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    RECT 0.27 -0.09 0.45 0.09 ;
END M10_M9_2x1_HV_E

VIA M10_M9_2x1_HV_W DEFAULT
  LAYER Metal9 ;
    RECT -0.49 -0.105 0.13 0.105 ;
  LAYER Metal10 ;
    RECT -0.48 -0.14 0.12 0.14 ;
  LAYER Via9 ;
    RECT -0.45 -0.09 -0.27 0.09 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_2x1_HV_W

VIA M10_M9_1x2_HV_N DEFAULT
  LAYER Metal9 ;
    RECT -0.13 -0.105 0.13 0.465 ;
  LAYER Metal10 ;
    RECT -0.12 -0.14 0.12 0.5 ;
  LAYER Via9 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    RECT -0.09 0.27 0.09 0.45 ;
END M10_M9_1x2_HV_N

VIA M10_M9_1x2_HV_S DEFAULT
  LAYER Metal9 ;
    RECT -0.13 -0.465 0.13 0.105 ;
  LAYER Metal10 ;
    RECT -0.12 -0.5 0.12 0.14 ;
  LAYER Via9 ;
    RECT -0.09 -0.45 0.09 -0.27 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M10_M9_1x2_HV_S

VIA M11_M10_VH DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.13 0.105 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_VH

VIA M11_M10_HH DEFAULT
  LAYER Metal10 ;
    RECT -0.13 -0.105 0.13 0.105 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_HH

VIA M11_M10_HV DEFAULT
  LAYER Metal10 ;
    RECT -0.13 -0.105 0.13 0.105 ;
  LAYER Metal11 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_HV

VIA M11_M10_VV DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.13 0.105 0.13 ;
  LAYER Metal11 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_VV

VIA M11_M10_M_NH DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.13 0.105 0.35 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_M_NH

VIA M11_M10_M_SH DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.35 0.105 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_M_SH

VIA M11_M10_2x1_VH_E DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.13 0.465 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.5 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    RECT 0.27 -0.09 0.45 0.09 ;
END M11_M10_2x1_VH_E

VIA M11_M10_2x1_VH_W DEFAULT
  LAYER Metal10 ;
    RECT -0.465 -0.13 0.105 0.13 ;
  LAYER Metal11 ;
    RECT -0.5 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.45 -0.09 -0.27 0.09 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_2x1_VH_W

VIA M11_M10_1x2_VH_N DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.13 0.105 0.49 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.48 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    RECT -0.09 0.27 0.09 0.45 ;
END M11_M10_1x2_VH_N

VIA M11_M10_1x2_VH_S DEFAULT
  LAYER Metal10 ;
    RECT -0.105 -0.49 0.105 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.48 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.45 0.09 -0.27 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_1x2_VH_S

VIA M2_M1_2x1_HH_E DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.04 0.23 0.04 ;
  LAYER Metal2 ;
    RECT -0.04 -0.04 0.23 0.04 ;
  LAYER Via1 ;
    RECT -0.01 -0.035 0.06 0.035 ;
    RECT 0.13 -0.035 0.2 0.035 ;
END M2_M1_2x1_HH_E

VIA M2_M1_2x1_HH_W DEFAULT
  LAYER Metal1 ;
    RECT -0.23 -0.04 0.04 0.04 ;
  LAYER Metal2 ;
    RECT -0.23 -0.04 0.04 0.04 ;
  LAYER Via1 ;
    RECT -0.2 -0.035 -0.13 0.035 ;
    RECT -0.06 -0.035 0.01 0.035 ;
END M2_M1_2x1_HH_W

VIA M2_M1_2x1_HH_C DEFAULT
  LAYER Metal1 ;
    RECT -0.135 -0.04 0.135 0.04 ;
  LAYER Metal2 ;
    RECT -0.135 -0.04 0.135 0.04 ;
  LAYER Via1 ;
    RECT -0.105 -0.035 -0.035 0.035 ;
    RECT 0.035 -0.035 0.105 0.035 ;
END M2_M1_2x1_HH_C

VIA M2_M1_1x2_VV_N DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.04 0.04 0.23 ;
  LAYER Metal2 ;
    RECT -0.04 -0.04 0.04 0.23 ;
  LAYER Via1 ;
    RECT -0.035 -0.01 0.035 0.06 ;
    RECT -0.035 0.13 0.035 0.2 ;
END M2_M1_1x2_VV_N

VIA M2_M1_1x2_VV_S DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.23 0.04 0.04 ;
  LAYER Metal2 ;
    RECT -0.04 -0.23 0.04 0.04 ;
  LAYER Via1 ;
    RECT -0.035 -0.2 0.035 -0.13 ;
    RECT -0.035 -0.06 0.035 0.01 ;
END M2_M1_1x2_VV_S

VIA M2_M1_1x2_VV_C DEFAULT
  LAYER Metal1 ;
    RECT -0.04 -0.135 0.04 0.135 ;
  LAYER Metal2 ;
    RECT -0.04 -0.135 0.04 0.135 ;
  LAYER Via1 ;
    RECT -0.035 -0.105 0.035 -0.035 ;
    RECT -0.035 0.035 0.035 0.105 ;
END M2_M1_1x2_VV_C

VIA M2_M1_2x2_HV DEFAULT
  LAYER Metal1 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Metal2 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Via1 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M2_M1_2x2_HV

VIA M3_M2_2x2_VH DEFAULT
  LAYER Metal2 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Metal3 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Via2 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M3_M2_2x2_VH

VIA M4_M3_2x2_HV DEFAULT
  LAYER Metal3 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Metal4 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Via3 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M4_M3_2x2_HV

VIA M5_M4_2x2_VH DEFAULT
  LAYER Metal4 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Metal5 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Via4 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M5_M4_2x2_VH

VIA M6_M5_2x2_HV DEFAULT
  LAYER Metal5 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Metal6 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Via5 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M6_M5_2x2_HV

VIA M7_M6_2x2_VH DEFAULT
  LAYER Metal6 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Metal7 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Via6 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M7_M6_2x2_VH

VIA M8_M7_2x2_HV DEFAULT
  LAYER Metal7 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Metal8 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Via7 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M8_M7_2x2_HV

VIA M9_M8_2x2_VH DEFAULT
  LAYER Metal8 ;
    RECT -0.125 -0.15 0.125 0.15 ;
  LAYER Metal9 ;
    RECT -0.15 -0.125 0.15 0.125 ;
  LAYER Via8 ;
    RECT -0.12 -0.12 -0.05 -0.05 ;
    RECT 0.05 -0.12 0.12 -0.05 ;
    RECT -0.12 0.05 -0.05 0.12 ;
    RECT 0.05 0.05 0.12 0.12 ;
END M9_M8_2x2_VH

VIA M10_M9_2x2_HV DEFAULT
  LAYER Metal9 ;
    RECT -0.32 -0.295 0.32 0.295 ;
  LAYER Metal10 ;
    RECT -0.31 -0.33 0.31 0.33 ;
  LAYER Via9 ;
    RECT -0.28 -0.28 -0.1 -0.1 ;
    RECT 0.1 -0.28 0.28 -0.1 ;
    RECT -0.28 0.1 -0.1 0.28 ;
    RECT 0.1 0.1 0.28 0.28 ;
END M10_M9_2x2_HV

VIA M11_M10_VH_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.13 0.11 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_VH_NEW

VIA M11_M10_HH_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.13 -0.11 0.13 0.11 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_HH_NEW

VIA M11_M10_HV_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.13 -0.11 0.13 0.11 ;
  LAYER Metal11 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_HV_NEW

VIA M11_M10_VV_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.13 0.11 0.13 ;
  LAYER Metal11 ;
    RECT -0.12 -0.14 0.12 0.14 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_VV_NEW

VIA M11_M10_M_NH_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.13 0.11 0.33 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_M_NH_NEW

VIA M11_M10_M_SH_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.33 0.11 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_M_SH_NEW

VIA M11_M10_1x2_VH_N_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.13 0.11 0.49 ;
  LAYER Metal11 ;
    RECT -0.14 -0.12 0.14 0.48 ;
  LAYER Via10 ;
    RECT -0.09 -0.09 0.09 0.09 ;
    RECT -0.09 0.27 0.09 0.45 ;
END M11_M10_1x2_VH_N_NEW

VIA M11_M10_1x2_VH_S_NEW DEFAULT
  LAYER Metal10 ;
    RECT -0.11 -0.49 0.11 0.13 ;
  LAYER Metal11 ;
    RECT -0.14 -0.48 0.14 0.12 ;
  LAYER Via10 ;
    RECT -0.09 -0.45 0.09 -0.27 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M11_M10_1x2_VH_S_NEW

NONDEFAULTRULE LEFSpecialRouteSpec
  LAYER Metal1
    WIDTH 0.06 ;
  END Metal1
  LAYER Metal2
    WIDTH 0.08 ;
  END Metal2
  LAYER Metal3
    WIDTH 0.08 ;
  END Metal3
  LAYER Metal4
    WIDTH 0.08 ;
  END Metal4
  LAYER Metal5
    WIDTH 0.08 ;
  END Metal5
  LAYER Metal6
    WIDTH 0.08 ;
  END Metal6
  LAYER Metal7
    WIDTH 0.08 ;
  END Metal7
  LAYER Metal8
    WIDTH 0.08 ;
  END Metal8
  LAYER Metal9
    WIDTH 0.08 ;
  END Metal9
  LAYER Metal10
    WIDTH 0.22 ;
  END Metal10
  LAYER Metal11
    WIDTH 0.22 ;
  END Metal11
  USEVIARULE M2_M1 ;
  USEVIARULE M3_M2 ;
  USEVIARULE M4_M3 ;
  USEVIARULE M5_M4 ;
  USEVIARULE M6_M5 ;
  USEVIARULE M7_M6 ;
  USEVIARULE M8_M7 ;
  USEVIARULE M9_M8 ;
  USEVIARULE M10_M9 ;
  USEVIARULE M11_M10 ;
END LEFSpecialRouteSpec
NONDEFAULTRULE VLMDefaultSetup
  LAYER Metal1
    WIDTH 0.06 ;
  END Metal1
  LAYER Metal2
    WIDTH 0.08 ;
  END Metal2
  LAYER Metal3
    WIDTH 0.08 ;
  END Metal3
  LAYER Metal4
    WIDTH 0.08 ;
  END Metal4
  LAYER Metal5
    WIDTH 0.08 ;
  END Metal5
  LAYER Metal6
    WIDTH 0.08 ;
  END Metal6
  LAYER Metal7
    WIDTH 0.08 ;
  END Metal7
  LAYER Metal8
    WIDTH 0.08 ;
  END Metal8
  LAYER Metal9
    WIDTH 0.08 ;
  END Metal9
  LAYER Metal10
    WIDTH 0.22 ;
  END Metal10
  LAYER Metal11
    WIDTH 0.22 ;
  END Metal11
  USEVIARULE M1_PO ;
  USEVIARULE M1_NWELL ;
  USEVIARULE M1_PSUB ;
  USEVIARULE M1_NIMP ;
  USEVIARULE M1_PIMP ;
  USEVIARULE M1_DIFF ;
  USEVIARULE M2_M1 ;
  USEVIARULE M3_M2 ;
  USEVIARULE M4_M3 ;
  USEVIARULE M5_M4 ;
  USEVIARULE M6_M5 ;
  USEVIARULE M7_M6 ;
  USEVIARULE M8_M7 ;
  USEVIARULE M9_M8 ;
  USEVIARULE M10_M9 ;
  USEVIARULE M11_M10 ;
END VLMDefaultSetup
SITE CoreSite
  CLASS CORE ;
  SIZE 0.2 BY 1.71 ;
END CoreSite

SITE IOSite
  CLASS PAD ;
  SIZE 1 BY 240 ;
END IOSite

SITE CornerSite
  CLASS PAD ;
  SIZE 240 BY 240 ;
END CornerSite

SITE CoreSiteDouble
  CLASS CORE ;
  SIZE 0.2 BY 3.42 ;
END CoreSiteDouble

END LIBRARY
